`timescale 1ns/1ns

/*
MIPI CSI RX to Parallel Bridge (c) by Gaurav Singh www.CircuitValley.com

MIPI CSI RX to Parallel Bridge is licensed under a
Creative Commons Attribution 3.0 Unported License.

You should have received a copy of the license along with this
work.  If not, see <http://creativecommons.org/licenses/by/3.0/>.
*/

/*
Takes 64bit 4pixel yuv input from rgb2yuv module @ mipi byte clock outputs 32bit 2pixel yuv output @output_clk_i , 
output_clk_i must be generated by same way as mipi byte clock, output_clk_i must be exactly double to mipi byteclock
This implementation of Output reformatter outputs data which which meant to send out of the system to a 32bit receiver 
depending on requirement this will be need to be adapted as per the receiver 
*/

module output_reformatter(clk_i, //data changes on negedge 
						  output_clk_i, //output clock double to clk_i to get in 64bit and output 32bit
						  data_i,
						  data_in_valid_i,
						  output_o,
						  output_valid_o
						  );
						  

input clk_i;
input data_in_valid_i;
input [63:0]data_i;
output reg output_valid_o;
output reg [31:0]output_o;
input output_clk_i;

reg lsw; //select if lower 32bit or higher 32bit 

always @(posedge output_clk_i)
begin
	if (!data_in_valid_i)
	begin
		lsw <= 1'd0;
		output_valid_o <= 1'd0;
	end
	else
	begin
		lsw <= !lsw;
		output_valid_o <= 1'd1;
		output_o <= data_i[((lsw)?6'd0:6'd32) +:32];
	end
end

endmodule